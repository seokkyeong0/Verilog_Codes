// Code your design here
`include "Downscaler.sv"
`include "DS_Gray.sv"
`include "DS_Bypass.sv"
`include "DS_Sampling.sv"
`include "DS_Average.sv"
`include "DS_Average_3x3.sv"
`include "DS_Cross.sv"